library verilog;
use verilog.vl_types.all;
entity sti is
end sti;
