module sti_test;
  
  reg [9:0]in;
  reg [2:0]a1,a2;
  reg clk,reset;
  wire [39:0]out;
  
  initial
  begin
	clk <= 1;
	reset <= 0;
	a1 <= 3'b001;
	a2 <= 3'b111;
	#20
	reset <= 1;
	//#30
  in <= 10'b0000111101;
  end

  always #5 clk <= ~clk;

  test TEST1(in,out,a1,a2,clk,reset); // define input & output ports of your top module by youself 



endmodule