library verilog;
use verilog.vl_types.all;
entity sti_version is
end sti_version;
