library verilog;
use verilog.vl_types.all;
entity sti_decoding is
end sti_decoding;
