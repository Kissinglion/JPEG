library verilog;
use verilog.vl_types.all;
entity sti_zig is
end sti_zig;
