library verilog;
use verilog.vl_types.all;
entity sti_test is
end sti_test;
