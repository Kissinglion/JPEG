module RLE2();
  
  input [63:0]in;
  output
  
  wire [223:0]out_temp;
  
  always@(*)
  begin
    if(next==0)
      
  
  
  
  assign out = {count,a[i]};
  
  assign out_temp = out_temp<<i + out;
  
  
  //SRAM512x16 MEM_OUT(1'b0,out_temp[111:0],11'd0,count3[3:0]-4'b0010,1'b0,clk, DO);