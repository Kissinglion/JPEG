library verilog;
use verilog.vl_types.all;
entity sti_project2 is
end sti_project2;
