library verilog;
use verilog.vl_types.all;
entity top_memory_test is
    port(
        clk             : in     vl_logic;
        reset           : in     vl_logic
    );
end top_memory_test;
