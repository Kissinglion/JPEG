library verilog;
use verilog.vl_types.all;
entity sti_rle2 is
end sti_rle2;
