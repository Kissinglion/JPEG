module sti;


reg clk;
reg reset;
reg [79:0]in;
wire [319:0]out;
//wire [2:0]run;

initial
begin
	clk <= 1;
	reset <= 0;
	#20
	reset <= 1;
	//#30
  in <= 80'h42_01_00_00_00_00_00_00_00_00;
  #10
  in <= 80'h00_00_00_00_00_00_0C_00_00_00;
  #10
  in <= 80'h00_00_00_00_00_00_00_00_00_00;
  #10
  in <= 80'h0B_FF_00_00_00_00_00_00_00_00;
  #10
  in <= 80'h01_FF_00_DD_00_00_00_00_00_00;
  #10
  in <= 80'h00_00_01_DD_00_00_00_00_00_00;
  #10
  in <= 80'h00_00_07_00_00_00_00_00_00_00;
  #10
  in <= 80'h00_00_00_00_00_00_00_00_00_00;
  //stage2
  
  #10
  in <= 64'h42_04_00_00_0D_00_00_00;
  #10
  in <= 64'h00_0C_00_03_00_00_00_00;
  #10
  in <= 64'hF2_00_00_00_00_00_07_00;
  #10
  in <= 64'h0B_FF_00_00_00_00_00_00;
  #10
  in <= 64'h01_FF_00_00_00_00_00_00;
  #10
  in <= 64'h00_00_00_00_00_00_00_00;
  #10
  in <= 64'h00_00_00_00_00_00_00_07;
  #10
  in <= 64'h00_00_00_00_00_00_00_00;
  
end

always #5 clk <= ~clk;

RLE_top TEST(in,out,clk,reset); // define input & output ports of your top module by youself 



endmodule

