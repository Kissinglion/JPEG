library verilog;
use verilog.vl_types.all;
entity sti_quant is
end sti_quant;
