module top_memory_test (clk,reset);
  
  input clk,reset;

  
  wire [15:0]count1;
  wire [14:0]count2,count3;
<<<<<<< HEAD

  wire [71:0]DCT_out1,tp_out1,tp_out2;
  wire [79:0]DCT_out2,DCT_out2_ff;
  wire [63:0]DIN1;
	wire [71:0]DIN2;
  wire [63:0]qt_out,DO,tp_out4,tp_out3,out;
  wire [111:0]rle_out;
  wire en1,en2,en3,en_rle;
=======
  wire [71:0]DCT_out1,tp_out1,tp_out2,DIN2;
  wire [79:0]DCT_out2,DO1,out1,DCT_out2_ff;
  wire [63:0]DIN1;
  wire [63:0]qt_out,qt_out1,zg_out1,zg_out2,zg_out,DO,tp_out3,tp_out4,out;
  wire en1,en2,en3;
>>>>>>> 08994d5726a6be19c6546bf350c9c3cf88d5c7a4
  wire [191:0]out_temp;
  wire [111:0]rle_out,rle_out1;
  wire en_rle;
  wire [79:0]tp_out33,tp_out44;

  
  SRAM32768x64 MEM_IN(1'b1,64'b0,count1[14:4],count1[3:0],1'b0,clk, DIN1 );
  
  DCT_first     d1(DIN1,DCT_out1);
  
  //D_ff_80b      d3(DCT_out2,DCT_out2_ff,clk,reset);
  
  Quantization_re qt(DCT_out2,qt_out,(count1[2:0]-3'b010),clk,reset);
  
  TPmem1 TP1(DCT_out1, en1,clk,reset,tp_out1);
  TPmem1 TP2(DCT_out1,~en1,clk,reset,tp_out2);
<<<<<<< HEAD

	DCT_second    d2(DIN2,DCT_out2,count1[2:0]);

	D_ff_80b				df1(DCT_out2,DCT_out2_ff,clk,reset);
	Quantization_re qt2(DCT_out2_ff,qt_out,(count1[2:0]-3'b011),clk,reset);

	ZigZag_TP	Zg3(qt_out, en2,clk,reset,tp_out3),
						Zg4(qt_out,~en2,clk,reset,tp_out4);

	SRAM32768x64 MEM_OUT(1'b0,out,count2[14:4],count2[3:0],1'b0,clk, DO);

  RLE_top  rl(out,rle_out,clk,en_rle);   
=======
  
  ZigZag_TP TP3(qt_out,  en2,clk,reset,tp_out3),
            TP4(qt_out, ~en2,clk,reset,tp_out4);
  
           
  RLE_top3  rl(out,rle_out,clk,en_rle);         
  
           
  TPmem2 TP5(DCT_out2, en2,clk,reset,tp_out33);
  TPmem2 TP6(DCT_out2,~en2,clk,reset,tp_out44);
  
  ZigZag  Zg1(qt_out1, en3,clk,reset,zg_out1);
  ZigZag  Zg2(qt_out1,~en3,clk,reset,zg_out2);
  
  Quantization qt1(out1,qt_out1,(count1[2:0]-3'b011),clk,reset);
  
  RLE_top3  rl1(zg_out,rle_out1,clk,en_rle1);
  
>>>>>>> 08994d5726a6be19c6546bf350c9c3cf88d5c7a4
  
  counter  cnt1(count1,       clk,reset);
  counter2 cnt2(count1,count2,clk,reset);
  counter3 cnt3(count1,count3,clk,reset);
  
  TPcontrol tp1(count1[4:0],en1,en2,en3,clk,reset);
  
<<<<<<< HEAD
  assign en_rle = (count1>=19)? 1'b1 : 1'b0;
  assign DIN2 = en1 ? tp_out2 : tp_out1;
	assign out = en2 ? tp_out4 : tp_out3;
=======
  
  
  assign en_rle = (count1>=18)? 1'b1 : 1'b0;
  assign en_rle1 = (count1>=27)? 1'b1 : 1'b0;
  assign DIN2 = en1 ? tp_out2 : tp_out1;
  assign out =  en2 ? tp_out4 : tp_out3;
  assign out1 = en2 ? tp_out44 : tp_out33;
  assign zg_out = en3 ? zg_out2 : zg_out1;
>>>>>>> 08994d5726a6be19c6546bf350c9c3cf88d5c7a4
endmodule

module counter(count,clk,reset);
  
  input clk,reset;
  output reg [15:0]count;
  
  always @(posedge clk)
  begin
    if(~reset)
      count <= 16'b0;
    else
      if(count == 16'b1111111111111111)
        count <= count;
      else
        count <= count + 1'b1;
  end
endmodule

module counter2(count1,count2,clk,reset);
  
  input clk,reset;
  input [15:0]count1;
  output reg [14:0]count2;
  
  always @(posedge clk)
  begin
    if(~reset)
      count2 <= 15'b0;
    else
      begin
        if(count1 <= 16'h0013)//27
          count2 <= 15'b0;
        else
          begin
            if(count2 == 15'b111111111111111)
              count2 <= count2;
            else
              count2 <= count2 + 1'b1;
          end
      end
  end
endmodule

module counter3(count1,count2,clk,reset);
  
  input clk,reset;
  input [15:0]count1;
  output reg [14:0]count2;
  
  always @(posedge clk)
  begin
    if(~reset)
      count2 <= 15'b0;
    else
      begin
        if(count1 <= 16'h0012)//18
          count2 <= 15'b0;
        else
          begin
            if(count2 == 15'b111111111111111)
              count2 <= count2;
            else
              count2 <= count2 + 1'b1;
          end
      end
  end
endmodule
     
module TPcontrol(count,en1,en2,en3,clk,reset);
  
input [4:0]count;
input clk,reset;
output reg en1,en2,en3;
  
  always @(posedge clk)
  begin
    if(count[3:0] == 4'b0000)
      en1 <= 1'b1;
    else
      begin
        if(count[2:0] == 3'b000)      
          en1 <= ~en1;
      end
  end

  always @(posedge clk)
    if(count[3:0]==4'b1010)
      	en2<=1'b1;
    else if(count[2:0] == 3'b010)
        en2<=(~en2);
        
  always @(posedge clk)
  begin
    if (count == 5'b10010)
      en3 <=1'b1;
    else if (count[2:0] == 3'b010)
      en3 <= (~en3);
  end
    
endmodule